`timescale 1ns/1ns

module testbench();

    initial begin
        $finish();
    end

endmodule
