module z1top();

endmodule
