module z1top(
    input sysclk,
    output PMOD_CS,
    output PMOD_MOSI,
    output PMOD_SCK,
    output PMOD_DC,
    output PMOD_RES,
    output PMOD_VCCEN,
    output PMOD_EN
);

endmodule
